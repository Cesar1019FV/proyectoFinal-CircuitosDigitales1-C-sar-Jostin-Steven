`timescale 1ns / 1ps

module celda_final(
    input f_mid,
    output f
);

assign f = f_mid;

endmodule