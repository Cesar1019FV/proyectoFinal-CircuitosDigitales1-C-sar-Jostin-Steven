module CeldaFinalBit(output Z_out,
input P_mid
);

    not not_gate(Z_out, P_mid);

endmodule
